module counter(reset, gray, clock, out);

    input reset, gray, clock; // تعریف ورودی‌ها: reset, gray, و clock
    output reg [3:0] out; // تعریف خروجی out به عنوان یک رجیستر 4 بیتی
    reg [3:0] q; // تعریف یک رجیستر داخلی 4 بیتی به نام q

    // بلاک always که با لبه مثبت کلاک فعال می‌شود
    always @(posedge clock) begin
        if (reset) begin
            q <= 4'b0000; // اگر سیگنال reset فعال باشد، q را به 0 می‌بریم
        end else if (gray) begin
            // بخشی برای پیاده‌سازی کانتر گری کد
            case(q)
                // هر کیس، مقدار بعدی q را بر اساس الگوی گری کد تعیین می‌کند
                4'b0000: q <= 4'b0001;
                4'b0001: q <= 4'b0011;
                4'b0011: q <= 4'b0010;
                4'b0010: q <= 4'b0110;
                4'b0110: q <= 4'b0111;
                4'b0111: q <= 4'b0101;
                4'b0101: q <= 4'b0100;
                4'b0100: q <= 4'b1100;
                4'b1100: q <= 4'b1101;
                4'b1101: q <= 4'b1111;
                4'b1111: q <= 4'b1110;
                4'b1110: q <= 4'b1010;
                4'b1010: q <= 4'b1011;
                4'b1011: q <= 4'b1001;
                4'b1001: q <= 4'b1000;
                4'b1000: q <= 4'b0000;
                default: q <= 4'b0000; // در صورتی که مقدار q خارج از محدوده باشد، به صفر ریست می‌شود
            endcase
        end else begin
                // بخشی برای افزایش q در صورتی که gray فعال نباشد
                if (q == 4'b1111) begin
                    q <= 4'b0000; // اگر q به مقدار حداکثر رسیده باشد، به صفر برمی‌گردد
                end else 
                    q <= q + 1; // در غیر این صورت، q را یک واحد افزایش می‌دهیم
                
        end

        // انتقال مقدار q به خروجی out
    	assign out = q; // این خط، مقدار فعلی q را به خروجی out منتقل می‌کند
    end

endmodule